// Peripheral parameters
`define SPI_INST_NUM     2
`define SPI_NUM_CS       4
`define I2C_INST_NUM     2
`define PWM_INST_NUM     4
`define TIM_INST_NUM     4
`define UART_INST_NUM    4
`define SD_INST_NUM      4
`define QEM_INST_NUM     4
`define NUM_PINS        24
`define NUM_SPI_REGS     5
`define NUM_I2C_REGS     6
`define NUM_PWM_REGS     4
`define NUM_TIM_REGS     6
`define NUM_UART_REGS    6
`define NUM_SD_REGS     10
`define NUM_QEM_REGS     6
`define SPI_NUM_INTER    1
`define I2C_NUM_INTER    1
`define TIM_NUM_INTER    1
`define UART_NUM_INTER   2
`define SD_NUM_INTER     1
`define QEM_NUM_INTER    2
`define GPIO_NUM_INTER   1
`define NUM_INTER       52

// GPIO Config bit fields
`define MOD1_POS         9
`define MOD0_POS         8
`define SEL1_POS         7
`define SEL0_POS         6
`define IRQEN_POS        5
`define IRQPOL_POS       4
`define INTR_POS         3
`define IRQRES_POS       2
`define DATA_IN_POS      1
`define DATA_OUT_POS     0
