magic
tech sky130A
magscale 1 2
timestamp 1699253876
<< obsli1 >>
rect 1104 2159 582820 701777
<< obsm1 >>
rect 382 1504 583450 701956
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 110 703464 8030 703520
rect 8254 703464 24222 703520
rect 24446 703464 40414 703520
rect 40638 703464 56698 703520
rect 56922 703464 72890 703520
rect 73114 703464 89082 703520
rect 89306 703464 105366 703520
rect 105590 703464 121558 703520
rect 121782 703464 137750 703520
rect 137974 703464 154034 703520
rect 154258 703464 170226 703520
rect 170450 703464 186418 703520
rect 186642 703464 202702 703520
rect 202926 703464 218894 703520
rect 219118 703464 235086 703520
rect 235310 703464 251370 703520
rect 251594 703464 267562 703520
rect 267786 703464 283754 703520
rect 283978 703464 300038 703520
rect 300262 703464 316230 703520
rect 316454 703464 332422 703520
rect 332646 703464 348706 703520
rect 348930 703464 364898 703520
rect 365122 703464 381090 703520
rect 381314 703464 397374 703520
rect 397598 703464 413566 703520
rect 413790 703464 429758 703520
rect 429982 703464 446042 703520
rect 446266 703464 462234 703520
rect 462458 703464 478426 703520
rect 478650 703464 494710 703520
rect 494934 703464 510902 703520
rect 511126 703464 527094 703520
rect 527318 703464 543378 703520
rect 543602 703464 559570 703520
rect 559794 703464 575762 703520
rect 575986 703464 583444 703520
rect 110 536 583444 703464
rect 110 54 486 536
rect 710 54 1590 536
rect 1814 54 2786 536
rect 3010 54 3982 536
rect 4206 54 5178 536
rect 5402 54 6374 536
rect 6598 54 7570 536
rect 7794 54 8674 536
rect 8898 54 9870 536
rect 10094 54 11066 536
rect 11290 54 12262 536
rect 12486 54 13458 536
rect 13682 54 14654 536
rect 14878 54 15850 536
rect 16074 54 16954 536
rect 17178 54 18150 536
rect 18374 54 19346 536
rect 19570 54 20542 536
rect 20766 54 21738 536
rect 21962 54 22934 536
rect 23158 54 24130 536
rect 24354 54 25234 536
rect 25458 54 26430 536
rect 26654 54 27626 536
rect 27850 54 28822 536
rect 29046 54 30018 536
rect 30242 54 31214 536
rect 31438 54 32318 536
rect 32542 54 33514 536
rect 33738 54 34710 536
rect 34934 54 35906 536
rect 36130 54 37102 536
rect 37326 54 38298 536
rect 38522 54 39494 536
rect 39718 54 40598 536
rect 40822 54 41794 536
rect 42018 54 42990 536
rect 43214 54 44186 536
rect 44410 54 45382 536
rect 45606 54 46578 536
rect 46802 54 47774 536
rect 47998 54 48878 536
rect 49102 54 50074 536
rect 50298 54 51270 536
rect 51494 54 52466 536
rect 52690 54 53662 536
rect 53886 54 54858 536
rect 55082 54 55962 536
rect 56186 54 57158 536
rect 57382 54 58354 536
rect 58578 54 59550 536
rect 59774 54 60746 536
rect 60970 54 61942 536
rect 62166 54 63138 536
rect 63362 54 64242 536
rect 64466 54 65438 536
rect 65662 54 66634 536
rect 66858 54 67830 536
rect 68054 54 69026 536
rect 69250 54 70222 536
rect 70446 54 71418 536
rect 71642 54 72522 536
rect 72746 54 73718 536
rect 73942 54 74914 536
rect 75138 54 76110 536
rect 76334 54 77306 536
rect 77530 54 78502 536
rect 78726 54 79606 536
rect 79830 54 80802 536
rect 81026 54 81998 536
rect 82222 54 83194 536
rect 83418 54 84390 536
rect 84614 54 85586 536
rect 85810 54 86782 536
rect 87006 54 87886 536
rect 88110 54 89082 536
rect 89306 54 90278 536
rect 90502 54 91474 536
rect 91698 54 92670 536
rect 92894 54 93866 536
rect 94090 54 95062 536
rect 95286 54 96166 536
rect 96390 54 97362 536
rect 97586 54 98558 536
rect 98782 54 99754 536
rect 99978 54 100950 536
rect 101174 54 102146 536
rect 102370 54 103250 536
rect 103474 54 104446 536
rect 104670 54 105642 536
rect 105866 54 106838 536
rect 107062 54 108034 536
rect 108258 54 109230 536
rect 109454 54 110426 536
rect 110650 54 111530 536
rect 111754 54 112726 536
rect 112950 54 113922 536
rect 114146 54 115118 536
rect 115342 54 116314 536
rect 116538 54 117510 536
rect 117734 54 118706 536
rect 118930 54 119810 536
rect 120034 54 121006 536
rect 121230 54 122202 536
rect 122426 54 123398 536
rect 123622 54 124594 536
rect 124818 54 125790 536
rect 126014 54 126894 536
rect 127118 54 128090 536
rect 128314 54 129286 536
rect 129510 54 130482 536
rect 130706 54 131678 536
rect 131902 54 132874 536
rect 133098 54 134070 536
rect 134294 54 135174 536
rect 135398 54 136370 536
rect 136594 54 137566 536
rect 137790 54 138762 536
rect 138986 54 139958 536
rect 140182 54 141154 536
rect 141378 54 142350 536
rect 142574 54 143454 536
rect 143678 54 144650 536
rect 144874 54 145846 536
rect 146070 54 147042 536
rect 147266 54 148238 536
rect 148462 54 149434 536
rect 149658 54 150538 536
rect 150762 54 151734 536
rect 151958 54 152930 536
rect 153154 54 154126 536
rect 154350 54 155322 536
rect 155546 54 156518 536
rect 156742 54 157714 536
rect 157938 54 158818 536
rect 159042 54 160014 536
rect 160238 54 161210 536
rect 161434 54 162406 536
rect 162630 54 163602 536
rect 163826 54 164798 536
rect 165022 54 165994 536
rect 166218 54 167098 536
rect 167322 54 168294 536
rect 168518 54 169490 536
rect 169714 54 170686 536
rect 170910 54 171882 536
rect 172106 54 173078 536
rect 173302 54 174182 536
rect 174406 54 175378 536
rect 175602 54 176574 536
rect 176798 54 177770 536
rect 177994 54 178966 536
rect 179190 54 180162 536
rect 180386 54 181358 536
rect 181582 54 182462 536
rect 182686 54 183658 536
rect 183882 54 184854 536
rect 185078 54 186050 536
rect 186274 54 187246 536
rect 187470 54 188442 536
rect 188666 54 189638 536
rect 189862 54 190742 536
rect 190966 54 191938 536
rect 192162 54 193134 536
rect 193358 54 194330 536
rect 194554 54 195526 536
rect 195750 54 196722 536
rect 196946 54 197826 536
rect 198050 54 199022 536
rect 199246 54 200218 536
rect 200442 54 201414 536
rect 201638 54 202610 536
rect 202834 54 203806 536
rect 204030 54 205002 536
rect 205226 54 206106 536
rect 206330 54 207302 536
rect 207526 54 208498 536
rect 208722 54 209694 536
rect 209918 54 210890 536
rect 211114 54 212086 536
rect 212310 54 213282 536
rect 213506 54 214386 536
rect 214610 54 215582 536
rect 215806 54 216778 536
rect 217002 54 217974 536
rect 218198 54 219170 536
rect 219394 54 220366 536
rect 220590 54 221470 536
rect 221694 54 222666 536
rect 222890 54 223862 536
rect 224086 54 225058 536
rect 225282 54 226254 536
rect 226478 54 227450 536
rect 227674 54 228646 536
rect 228870 54 229750 536
rect 229974 54 230946 536
rect 231170 54 232142 536
rect 232366 54 233338 536
rect 233562 54 234534 536
rect 234758 54 235730 536
rect 235954 54 236926 536
rect 237150 54 238030 536
rect 238254 54 239226 536
rect 239450 54 240422 536
rect 240646 54 241618 536
rect 241842 54 242814 536
rect 243038 54 244010 536
rect 244234 54 245114 536
rect 245338 54 246310 536
rect 246534 54 247506 536
rect 247730 54 248702 536
rect 248926 54 249898 536
rect 250122 54 251094 536
rect 251318 54 252290 536
rect 252514 54 253394 536
rect 253618 54 254590 536
rect 254814 54 255786 536
rect 256010 54 256982 536
rect 257206 54 258178 536
rect 258402 54 259374 536
rect 259598 54 260570 536
rect 260794 54 261674 536
rect 261898 54 262870 536
rect 263094 54 264066 536
rect 264290 54 265262 536
rect 265486 54 266458 536
rect 266682 54 267654 536
rect 267878 54 268758 536
rect 268982 54 269954 536
rect 270178 54 271150 536
rect 271374 54 272346 536
rect 272570 54 273542 536
rect 273766 54 274738 536
rect 274962 54 275934 536
rect 276158 54 277038 536
rect 277262 54 278234 536
rect 278458 54 279430 536
rect 279654 54 280626 536
rect 280850 54 281822 536
rect 282046 54 283018 536
rect 283242 54 284214 536
rect 284438 54 285318 536
rect 285542 54 286514 536
rect 286738 54 287710 536
rect 287934 54 288906 536
rect 289130 54 290102 536
rect 290326 54 291298 536
rect 291522 54 292494 536
rect 292718 54 293598 536
rect 293822 54 294794 536
rect 295018 54 295990 536
rect 296214 54 297186 536
rect 297410 54 298382 536
rect 298606 54 299578 536
rect 299802 54 300682 536
rect 300906 54 301878 536
rect 302102 54 303074 536
rect 303298 54 304270 536
rect 304494 54 305466 536
rect 305690 54 306662 536
rect 306886 54 307858 536
rect 308082 54 308962 536
rect 309186 54 310158 536
rect 310382 54 311354 536
rect 311578 54 312550 536
rect 312774 54 313746 536
rect 313970 54 314942 536
rect 315166 54 316138 536
rect 316362 54 317242 536
rect 317466 54 318438 536
rect 318662 54 319634 536
rect 319858 54 320830 536
rect 321054 54 322026 536
rect 322250 54 323222 536
rect 323446 54 324326 536
rect 324550 54 325522 536
rect 325746 54 326718 536
rect 326942 54 327914 536
rect 328138 54 329110 536
rect 329334 54 330306 536
rect 330530 54 331502 536
rect 331726 54 332606 536
rect 332830 54 333802 536
rect 334026 54 334998 536
rect 335222 54 336194 536
rect 336418 54 337390 536
rect 337614 54 338586 536
rect 338810 54 339782 536
rect 340006 54 340886 536
rect 341110 54 342082 536
rect 342306 54 343278 536
rect 343502 54 344474 536
rect 344698 54 345670 536
rect 345894 54 346866 536
rect 347090 54 347970 536
rect 348194 54 349166 536
rect 349390 54 350362 536
rect 350586 54 351558 536
rect 351782 54 352754 536
rect 352978 54 353950 536
rect 354174 54 355146 536
rect 355370 54 356250 536
rect 356474 54 357446 536
rect 357670 54 358642 536
rect 358866 54 359838 536
rect 360062 54 361034 536
rect 361258 54 362230 536
rect 362454 54 363426 536
rect 363650 54 364530 536
rect 364754 54 365726 536
rect 365950 54 366922 536
rect 367146 54 368118 536
rect 368342 54 369314 536
rect 369538 54 370510 536
rect 370734 54 371614 536
rect 371838 54 372810 536
rect 373034 54 374006 536
rect 374230 54 375202 536
rect 375426 54 376398 536
rect 376622 54 377594 536
rect 377818 54 378790 536
rect 379014 54 379894 536
rect 380118 54 381090 536
rect 381314 54 382286 536
rect 382510 54 383482 536
rect 383706 54 384678 536
rect 384902 54 385874 536
rect 386098 54 387070 536
rect 387294 54 388174 536
rect 388398 54 389370 536
rect 389594 54 390566 536
rect 390790 54 391762 536
rect 391986 54 392958 536
rect 393182 54 394154 536
rect 394378 54 395258 536
rect 395482 54 396454 536
rect 396678 54 397650 536
rect 397874 54 398846 536
rect 399070 54 400042 536
rect 400266 54 401238 536
rect 401462 54 402434 536
rect 402658 54 403538 536
rect 403762 54 404734 536
rect 404958 54 405930 536
rect 406154 54 407126 536
rect 407350 54 408322 536
rect 408546 54 409518 536
rect 409742 54 410714 536
rect 410938 54 411818 536
rect 412042 54 413014 536
rect 413238 54 414210 536
rect 414434 54 415406 536
rect 415630 54 416602 536
rect 416826 54 417798 536
rect 418022 54 418902 536
rect 419126 54 420098 536
rect 420322 54 421294 536
rect 421518 54 422490 536
rect 422714 54 423686 536
rect 423910 54 424882 536
rect 425106 54 426078 536
rect 426302 54 427182 536
rect 427406 54 428378 536
rect 428602 54 429574 536
rect 429798 54 430770 536
rect 430994 54 431966 536
rect 432190 54 433162 536
rect 433386 54 434358 536
rect 434582 54 435462 536
rect 435686 54 436658 536
rect 436882 54 437854 536
rect 438078 54 439050 536
rect 439274 54 440246 536
rect 440470 54 441442 536
rect 441666 54 442546 536
rect 442770 54 443742 536
rect 443966 54 444938 536
rect 445162 54 446134 536
rect 446358 54 447330 536
rect 447554 54 448526 536
rect 448750 54 449722 536
rect 449946 54 450826 536
rect 451050 54 452022 536
rect 452246 54 453218 536
rect 453442 54 454414 536
rect 454638 54 455610 536
rect 455834 54 456806 536
rect 457030 54 458002 536
rect 458226 54 459106 536
rect 459330 54 460302 536
rect 460526 54 461498 536
rect 461722 54 462694 536
rect 462918 54 463890 536
rect 464114 54 465086 536
rect 465310 54 466190 536
rect 466414 54 467386 536
rect 467610 54 468582 536
rect 468806 54 469778 536
rect 470002 54 470974 536
rect 471198 54 472170 536
rect 472394 54 473366 536
rect 473590 54 474470 536
rect 474694 54 475666 536
rect 475890 54 476862 536
rect 477086 54 478058 536
rect 478282 54 479254 536
rect 479478 54 480450 536
rect 480674 54 481646 536
rect 481870 54 482750 536
rect 482974 54 483946 536
rect 484170 54 485142 536
rect 485366 54 486338 536
rect 486562 54 487534 536
rect 487758 54 488730 536
rect 488954 54 489834 536
rect 490058 54 491030 536
rect 491254 54 492226 536
rect 492450 54 493422 536
rect 493646 54 494618 536
rect 494842 54 495814 536
rect 496038 54 497010 536
rect 497234 54 498114 536
rect 498338 54 499310 536
rect 499534 54 500506 536
rect 500730 54 501702 536
rect 501926 54 502898 536
rect 503122 54 504094 536
rect 504318 54 505290 536
rect 505514 54 506394 536
rect 506618 54 507590 536
rect 507814 54 508786 536
rect 509010 54 509982 536
rect 510206 54 511178 536
rect 511402 54 512374 536
rect 512598 54 513478 536
rect 513702 54 514674 536
rect 514898 54 515870 536
rect 516094 54 517066 536
rect 517290 54 518262 536
rect 518486 54 519458 536
rect 519682 54 520654 536
rect 520878 54 521758 536
rect 521982 54 522954 536
rect 523178 54 524150 536
rect 524374 54 525346 536
rect 525570 54 526542 536
rect 526766 54 527738 536
rect 527962 54 528934 536
rect 529158 54 530038 536
rect 530262 54 531234 536
rect 531458 54 532430 536
rect 532654 54 533626 536
rect 533850 54 534822 536
rect 535046 54 536018 536
rect 536242 54 537122 536
rect 537346 54 538318 536
rect 538542 54 539514 536
rect 539738 54 540710 536
rect 540934 54 541906 536
rect 542130 54 543102 536
rect 543326 54 544298 536
rect 544522 54 545402 536
rect 545626 54 546598 536
rect 546822 54 547794 536
rect 548018 54 548990 536
rect 549214 54 550186 536
rect 550410 54 551382 536
rect 551606 54 552578 536
rect 552802 54 553682 536
rect 553906 54 554878 536
rect 555102 54 556074 536
rect 556298 54 557270 536
rect 557494 54 558466 536
rect 558690 54 559662 536
rect 559886 54 560766 536
rect 560990 54 561962 536
rect 562186 54 563158 536
rect 563382 54 564354 536
rect 564578 54 565550 536
rect 565774 54 566746 536
rect 566970 54 567942 536
rect 568166 54 569046 536
rect 569270 54 570242 536
rect 570466 54 571438 536
rect 571662 54 572634 536
rect 572858 54 573830 536
rect 574054 54 575026 536
rect 575250 54 576222 536
rect 576446 54 577326 536
rect 577550 54 578522 536
rect 578746 54 579718 536
rect 579942 54 580914 536
rect 581138 54 582110 536
rect 582334 54 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 54 697540 583520 701997
rect 560 697404 583520 697540
rect 560 697140 583440 697404
rect 54 697004 583440 697140
rect 54 684484 583520 697004
rect 560 684084 583520 684484
rect 54 684076 583520 684084
rect 54 683676 583440 684076
rect 54 671428 583520 683676
rect 560 671028 583520 671428
rect 54 670884 583520 671028
rect 54 670484 583440 670884
rect 54 658372 583520 670484
rect 560 657972 583520 658372
rect 54 657556 583520 657972
rect 54 657156 583440 657556
rect 54 645316 583520 657156
rect 560 644916 583520 645316
rect 54 644228 583520 644916
rect 54 643828 583440 644228
rect 54 632260 583520 643828
rect 560 631860 583520 632260
rect 54 631036 583520 631860
rect 54 630636 583440 631036
rect 54 619340 583520 630636
rect 560 618940 583520 619340
rect 54 617708 583520 618940
rect 54 617308 583440 617708
rect 54 606284 583520 617308
rect 560 605884 583520 606284
rect 54 604380 583520 605884
rect 54 603980 583440 604380
rect 54 593228 583520 603980
rect 560 592828 583520 593228
rect 54 591188 583520 592828
rect 54 590788 583440 591188
rect 54 580172 583520 590788
rect 560 579772 583520 580172
rect 54 577860 583520 579772
rect 54 577460 583440 577860
rect 54 567116 583520 577460
rect 560 566716 583520 567116
rect 54 564532 583520 566716
rect 54 564132 583440 564532
rect 54 554060 583520 564132
rect 560 553660 583520 554060
rect 54 551340 583520 553660
rect 54 550940 583440 551340
rect 54 541004 583520 550940
rect 560 540604 583520 541004
rect 54 538012 583520 540604
rect 54 537612 583440 538012
rect 54 528084 583520 537612
rect 560 527684 583520 528084
rect 54 524684 583520 527684
rect 54 524284 583440 524684
rect 54 515028 583520 524284
rect 560 514628 583520 515028
rect 54 511492 583520 514628
rect 54 511092 583440 511492
rect 54 501972 583520 511092
rect 560 501572 583520 501972
rect 54 498164 583520 501572
rect 54 497764 583440 498164
rect 54 488916 583520 497764
rect 560 488516 583520 488916
rect 54 484836 583520 488516
rect 54 484436 583440 484836
rect 54 475860 583520 484436
rect 560 475460 583520 475860
rect 54 471644 583520 475460
rect 54 471244 583440 471644
rect 54 462804 583520 471244
rect 560 462404 583520 462804
rect 54 458316 583520 462404
rect 54 457916 583440 458316
rect 54 449748 583520 457916
rect 560 449348 583520 449748
rect 54 444988 583520 449348
rect 54 444588 583440 444988
rect 54 436828 583520 444588
rect 560 436428 583520 436828
rect 54 431796 583520 436428
rect 54 431396 583440 431796
rect 54 423772 583520 431396
rect 560 423372 583520 423772
rect 54 418468 583520 423372
rect 54 418068 583440 418468
rect 54 410716 583520 418068
rect 560 410316 583520 410716
rect 54 405140 583520 410316
rect 54 404740 583440 405140
rect 54 397660 583520 404740
rect 560 397260 583520 397660
rect 54 391948 583520 397260
rect 54 391548 583440 391948
rect 54 384604 583520 391548
rect 560 384204 583520 384604
rect 54 378620 583520 384204
rect 54 378220 583440 378620
rect 54 371548 583520 378220
rect 560 371148 583520 371548
rect 54 365292 583520 371148
rect 54 364892 583440 365292
rect 54 358628 583520 364892
rect 560 358228 583520 358628
rect 54 352100 583520 358228
rect 54 351700 583440 352100
rect 54 345572 583520 351700
rect 560 345172 583520 345572
rect 54 338772 583520 345172
rect 54 338372 583440 338772
rect 54 332516 583520 338372
rect 560 332116 583520 332516
rect 54 325444 583520 332116
rect 54 325044 583440 325444
rect 54 319460 583520 325044
rect 560 319060 583520 319460
rect 54 312252 583520 319060
rect 54 311852 583440 312252
rect 54 306404 583520 311852
rect 560 306004 583520 306404
rect 54 298924 583520 306004
rect 54 298524 583440 298924
rect 54 293348 583520 298524
rect 560 292948 583520 293348
rect 54 285596 583520 292948
rect 54 285196 583440 285596
rect 54 280292 583520 285196
rect 560 279892 583520 280292
rect 54 272404 583520 279892
rect 54 272004 583440 272404
rect 54 267372 583520 272004
rect 560 266972 583520 267372
rect 54 259076 583520 266972
rect 54 258676 583440 259076
rect 54 254316 583520 258676
rect 560 253916 583520 254316
rect 54 245748 583520 253916
rect 54 245348 583440 245748
rect 54 241260 583520 245348
rect 560 240860 583520 241260
rect 54 232556 583520 240860
rect 54 232156 583440 232556
rect 54 228204 583520 232156
rect 560 227804 583520 228204
rect 54 219228 583520 227804
rect 54 218828 583440 219228
rect 54 215148 583520 218828
rect 560 214748 583520 215148
rect 54 205900 583520 214748
rect 54 205500 583440 205900
rect 54 202092 583520 205500
rect 560 201692 583520 202092
rect 54 192708 583520 201692
rect 54 192308 583440 192708
rect 54 189036 583520 192308
rect 560 188636 583520 189036
rect 54 179380 583520 188636
rect 54 178980 583440 179380
rect 54 176116 583520 178980
rect 560 175716 583520 176116
rect 54 166052 583520 175716
rect 54 165652 583440 166052
rect 54 163060 583520 165652
rect 560 162660 583520 163060
rect 54 152860 583520 162660
rect 54 152460 583440 152860
rect 54 150004 583520 152460
rect 560 149604 583520 150004
rect 54 139532 583520 149604
rect 54 139132 583440 139532
rect 54 136948 583520 139132
rect 560 136548 583520 136948
rect 54 126204 583520 136548
rect 54 125804 583440 126204
rect 54 123892 583520 125804
rect 560 123492 583520 123892
rect 54 113012 583520 123492
rect 54 112612 583440 113012
rect 54 110836 583520 112612
rect 560 110436 583520 110836
rect 54 99684 583520 110436
rect 54 99284 583440 99684
rect 54 97780 583520 99284
rect 560 97380 583520 97780
rect 54 86356 583520 97380
rect 54 85956 583440 86356
rect 54 84860 583520 85956
rect 560 84460 583520 84860
rect 54 73164 583520 84460
rect 54 72764 583440 73164
rect 54 71804 583520 72764
rect 560 71404 583520 71804
rect 54 59836 583520 71404
rect 54 59436 583440 59836
rect 54 58748 583520 59436
rect 560 58348 583520 58748
rect 54 46508 583520 58348
rect 54 46108 583440 46508
rect 54 45692 583520 46108
rect 560 45292 583520 45692
rect 54 33316 583520 45292
rect 54 32916 583440 33316
rect 54 32636 583520 32916
rect 560 32236 583520 32636
rect 54 19988 583520 32236
rect 54 19588 583440 19988
rect 54 19580 583520 19588
rect 560 19180 583520 19580
rect 54 6796 583520 19180
rect 54 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 54 2143 583520 6260
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 1794 -7654 2414 711590
rect 5514 -7654 6134 711590
rect 9234 -7654 9854 711590
rect 12954 -7654 13574 711590
rect 16674 -7654 17294 711590
rect 20394 -7654 21014 711590
rect 24114 -7654 24734 711590
rect 27834 -7654 28454 711590
rect 37794 -7654 38414 711590
rect 41514 -7654 42134 711590
rect 45234 -7654 45854 711590
rect 48954 -7654 49574 711590
rect 52674 -7654 53294 711590
rect 56394 -7654 57014 711590
rect 60114 -7654 60734 711590
rect 63834 -7654 64454 711590
rect 73794 645956 74414 711590
rect 77514 645956 78134 711590
rect 81234 646140 81854 711590
rect 84954 645956 85574 711590
rect 88674 645956 89294 711590
rect 92394 646140 93014 711590
rect 96114 645956 96734 711590
rect 99834 645956 100454 711590
rect 109794 645956 110414 711590
rect 113514 646140 114134 711590
rect 117234 645956 117854 711590
rect 120954 646140 121574 711590
rect 124674 645956 125294 711590
rect 128394 646140 129014 711590
rect 132114 645956 132734 711590
rect 135834 646140 136454 711590
rect 145794 646140 146414 711590
rect 149514 645956 150134 711590
rect 153234 646140 153854 711590
rect 156954 645956 157574 711590
rect 160674 646140 161294 711590
rect 164394 645956 165014 711590
rect 168114 646140 168734 711590
rect 171834 645956 172454 711590
rect 181794 645956 182414 711590
rect 185514 645956 186134 711590
rect 189234 645956 189854 711590
rect 192954 645956 193574 711590
rect 196674 645956 197294 711590
rect 200394 645956 201014 711590
rect 204114 645956 204734 711590
rect 207834 645956 208454 711590
rect 73794 479058 74414 558736
rect 77514 479058 78134 558736
rect 81234 479058 81854 558736
rect 84954 479058 85574 558736
rect 88674 479242 89294 558552
rect 92394 479058 93014 558736
rect 96114 479058 96734 558736
rect 99834 479058 100454 558736
rect 109794 479058 110414 558736
rect 113514 479242 114134 558552
rect 117234 479058 117854 558736
rect 120954 479242 121574 558552
rect 124674 479058 125294 558736
rect 128394 479242 129014 558552
rect 132114 479058 132734 558736
rect 135834 479242 136454 558552
rect 145794 479242 146414 558552
rect 149514 479058 150134 558736
rect 153234 479242 153854 558552
rect 156954 479242 157574 558552
rect 160674 479242 161294 558552
rect 164394 479242 165014 558552
rect 168114 479242 168734 558552
rect 171834 479242 172454 558552
rect 181794 479242 182414 558552
rect 185514 479242 186134 558552
rect 189234 479058 189854 558736
rect 192954 479242 193574 558552
rect 196674 479058 197294 558736
rect 200394 479058 201014 558736
rect 204114 479058 204734 558736
rect 207834 479058 208454 558736
rect 73794 312164 74414 391838
rect 77514 312164 78134 391838
rect 81234 312348 81854 391654
rect 84954 312164 85574 391838
rect 88674 312164 89294 391838
rect 92394 312348 93014 391654
rect 96114 312164 96734 391838
rect 99834 312164 100454 391838
rect 109794 312164 110414 391838
rect 113514 312348 114134 391654
rect 117234 312164 117854 391838
rect 120954 312348 121574 391654
rect 124674 312164 125294 391838
rect 128394 312348 129014 391654
rect 132114 312164 132734 391838
rect 135834 312348 136454 391654
rect 145794 312348 146414 391654
rect 149514 312164 150134 391838
rect 153234 312348 153854 391654
rect 156954 312164 157574 391838
rect 160674 312348 161294 391654
rect 164394 312164 165014 391838
rect 168114 312348 168734 391654
rect 171834 312164 172454 391838
rect 181794 312164 182414 391838
rect 185514 312164 186134 391838
rect 189234 312164 189854 391838
rect 192954 312164 193574 391838
rect 196674 312164 197294 391838
rect 200394 312164 201014 391838
rect 204114 312164 204734 391838
rect 207834 312164 208454 391838
rect 73794 145264 74414 224944
rect 77514 145264 78134 224944
rect 81234 145264 81854 224944
rect 84954 145264 85574 224944
rect 88674 145448 89294 224760
rect 92394 145264 93014 224944
rect 96114 145264 96734 224944
rect 99834 145264 100454 224944
rect 109794 145264 110414 224944
rect 113514 145448 114134 224760
rect 117234 145264 117854 224944
rect 120954 145448 121574 224760
rect 124674 145264 125294 224944
rect 128394 145448 129014 224760
rect 132114 145264 132734 224944
rect 135834 145448 136454 224760
rect 145794 145448 146414 224760
rect 149514 145264 150134 224944
rect 153234 145448 153854 224760
rect 156954 145448 157574 224760
rect 160674 145448 161294 224760
rect 164394 145448 165014 224760
rect 168114 145448 168734 224760
rect 171834 145448 172454 224760
rect 181794 145448 182414 224760
rect 185514 145448 186134 224760
rect 189234 145264 189854 224944
rect 192954 145448 193574 224760
rect 196674 145264 197294 224944
rect 200394 145264 201014 224944
rect 204114 145264 204734 224944
rect 207834 145264 208454 224944
rect 73794 -7654 74414 58044
rect 77514 -7654 78134 58044
rect 81234 -7654 81854 57860
rect 84954 -7654 85574 58044
rect 88674 -7654 89294 58044
rect 92394 -7654 93014 58086
rect 96114 -7654 96734 58044
rect 99834 -7654 100454 58044
rect 109794 -7654 110414 58044
rect 113514 -7654 114134 57860
rect 117234 -7654 117854 58044
rect 120954 -7654 121574 57860
rect 124674 -7654 125294 58044
rect 128394 -7654 129014 57860
rect 132114 -7654 132734 58044
rect 135834 -7654 136454 57860
rect 145794 -7654 146414 57860
rect 149514 -7654 150134 58044
rect 153234 -7654 153854 57860
rect 156954 -7654 157574 58044
rect 160674 -7654 161294 57860
rect 164394 -7654 165014 58086
rect 168114 -7654 168734 57860
rect 171834 -7654 172454 58044
rect 181794 -7654 182414 58044
rect 185514 -7654 186134 58044
rect 189234 -7654 189854 58044
rect 192954 -7654 193574 58044
rect 196674 -7654 197294 58044
rect 200394 -7654 201014 58086
rect 204114 -7654 204734 58044
rect 207834 -7654 208454 58044
rect 217794 -7654 218414 711590
rect 221514 -7654 222134 711590
rect 225234 -7654 225854 711590
rect 228954 -7654 229574 711590
rect 232674 -7654 233294 711590
rect 236394 -7654 237014 711590
rect 240114 -7654 240734 711590
rect 243834 -7654 244454 711590
rect 253794 -7654 254414 711590
rect 257514 -7654 258134 711590
rect 261234 -7654 261854 711590
rect 264954 -7654 265574 711590
rect 268674 -7654 269294 711590
rect 272394 -7654 273014 711590
rect 276114 -7654 276734 711590
rect 279834 -7654 280454 711590
rect 289794 -7654 290414 711590
rect 293514 -7654 294134 711590
rect 297234 -7654 297854 711590
rect 300954 -7654 301574 711590
rect 304674 -7654 305294 711590
rect 308394 -7654 309014 711590
rect 312114 -7654 312734 711590
rect 315834 -7654 316454 711590
rect 325794 -7654 326414 711590
rect 329514 -7654 330134 711590
rect 333234 -7654 333854 711590
rect 336954 -7654 337574 711590
rect 340674 -7654 341294 711590
rect 344394 -7654 345014 711590
rect 348114 -7654 348734 711590
rect 351834 -7654 352454 711590
rect 361794 -7654 362414 711590
rect 365514 -7654 366134 711590
rect 369234 -7654 369854 711590
rect 372954 645956 373574 711590
rect 376674 645956 377294 711590
rect 380394 645956 381014 711590
rect 384114 645956 384734 711590
rect 387834 645956 388454 711590
rect 397794 645956 398414 711590
rect 401514 645956 402134 711590
rect 405234 646140 405854 711590
rect 408954 645956 409574 711590
rect 412674 646140 413294 711590
rect 416394 645956 417014 711590
rect 420114 646140 420734 711590
rect 423834 645956 424454 711590
rect 433794 645956 434414 711590
rect 437514 646140 438134 711590
rect 441234 645956 441854 711590
rect 444954 646140 445574 711590
rect 448674 645956 449294 711590
rect 452394 646140 453014 711590
rect 456114 645956 456734 711590
rect 459834 646140 460454 711590
rect 469794 646140 470414 711590
rect 473514 645956 474134 711590
rect 477234 645956 477854 711590
rect 480954 645956 481574 711590
rect 484674 645956 485294 711590
rect 488394 645956 489014 711590
rect 492114 645956 492734 711590
rect 495834 645956 496454 711590
rect 505794 645956 506414 711590
rect 509514 645956 510134 711590
rect 372954 479058 373574 558736
rect 376674 479058 377294 558736
rect 380394 479058 381014 558736
rect 384114 479058 384734 558736
rect 387834 479242 388454 558552
rect 397794 479242 398414 558552
rect 401514 479242 402134 558552
rect 405234 479242 405854 558552
rect 408954 479242 409574 558552
rect 412674 479242 413294 558552
rect 416394 479058 417014 558736
rect 420114 479242 420734 558552
rect 423834 479242 424454 558552
rect 433794 479058 434414 558736
rect 437514 479242 438134 558552
rect 441234 479058 441854 558736
rect 444954 479242 445574 558552
rect 448674 479058 449294 558736
rect 452394 479242 453014 558552
rect 456114 479058 456734 558736
rect 459834 479242 460454 558552
rect 469794 479242 470414 558552
rect 473514 479058 474134 558736
rect 477234 479242 477854 558552
rect 480954 479058 481574 558736
rect 484674 479058 485294 558736
rect 488394 479058 489014 558736
rect 492114 479058 492734 558736
rect 495834 479058 496454 558736
rect 505794 479058 506414 558736
rect 509514 479058 510134 558736
rect 372954 312164 373574 391838
rect 376674 312164 377294 391838
rect 380394 312164 381014 391838
rect 384114 312164 384734 391838
rect 387834 312164 388454 391838
rect 397794 312164 398414 391838
rect 401514 312164 402134 391838
rect 405234 312348 405854 391654
rect 408954 312164 409574 391838
rect 412674 312348 413294 391654
rect 416394 312164 417014 391838
rect 420114 312348 420734 391654
rect 423834 312164 424454 391838
rect 433794 312164 434414 391838
rect 437514 312348 438134 391654
rect 441234 312164 441854 391838
rect 444954 312348 445574 391654
rect 448674 312164 449294 391838
rect 452394 312348 453014 391654
rect 456114 312164 456734 391838
rect 459834 312348 460454 391654
rect 469794 312348 470414 391654
rect 473514 312164 474134 391838
rect 477234 312164 477854 391838
rect 480954 312164 481574 391838
rect 484674 312164 485294 391838
rect 488394 312164 489014 391838
rect 492114 312164 492734 391838
rect 495834 312164 496454 391838
rect 505794 312164 506414 391838
rect 509514 312164 510134 391838
rect 372954 145264 373574 224944
rect 376674 145264 377294 224944
rect 380394 145264 381014 224944
rect 384114 145264 384734 224944
rect 387834 145448 388454 224760
rect 397794 145448 398414 224760
rect 401514 145448 402134 224760
rect 405234 145448 405854 224760
rect 408954 145448 409574 224760
rect 412674 145448 413294 224760
rect 416394 145264 417014 224944
rect 420114 145448 420734 224760
rect 423834 145448 424454 224760
rect 433794 145264 434414 224944
rect 437514 145448 438134 224760
rect 441234 145264 441854 224944
rect 444954 145448 445574 224760
rect 448674 145264 449294 224944
rect 452394 145448 453014 224760
rect 456114 145264 456734 224944
rect 459834 145448 460454 224760
rect 469794 145448 470414 224760
rect 473514 145264 474134 224944
rect 477234 145448 477854 224760
rect 480954 145264 481574 224944
rect 484674 145264 485294 224944
rect 488394 145264 489014 224944
rect 492114 145264 492734 224944
rect 495834 145264 496454 224944
rect 505794 145264 506414 224944
rect 509514 145264 510134 224944
rect 372954 -7654 373574 58044
rect 376674 -7654 377294 58044
rect 380394 -7654 381014 58086
rect 384114 -7654 384734 58044
rect 387834 -7654 388454 58044
rect 397794 -7654 398414 58044
rect 401514 -7654 402134 58044
rect 405234 -7654 405854 57860
rect 408954 -7654 409574 58044
rect 412674 -7654 413294 57860
rect 416394 -7654 417014 58086
rect 420114 -7654 420734 57860
rect 423834 -7654 424454 58044
rect 433794 -7654 434414 58044
rect 437514 -7654 438134 57860
rect 441234 -7654 441854 58044
rect 444954 -7654 445574 57860
rect 448674 -7654 449294 58044
rect 452394 -7654 453014 57860
rect 456114 -7654 456734 58044
rect 459834 -7654 460454 57860
rect 469794 -7654 470414 57860
rect 473514 -7654 474134 58044
rect 477234 -7654 477854 58044
rect 480954 -7654 481574 58044
rect 484674 -7654 485294 58044
rect 488394 -7654 489014 58086
rect 492114 -7654 492734 58044
rect 495834 -7654 496454 58044
rect 505794 -7654 506414 58044
rect 509514 -7654 510134 58044
rect 513234 -7654 513854 711590
rect 516954 -7654 517574 711590
rect 520674 -7654 521294 711590
rect 524394 -7654 525014 711590
rect 528114 -7654 528734 711590
rect 531834 -7654 532454 711590
rect 541794 -7654 542414 711590
rect 545514 -7654 546134 711590
rect 549234 -7654 549854 711590
rect 552954 -7654 553574 711590
rect 556674 -7654 557294 711590
rect 560394 -7654 561014 711590
rect 564114 -7654 564734 711590
rect 567834 -7654 568454 711590
rect 577794 -7654 578414 711590
rect 581514 -7654 582134 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 59 2347 1714 701997
rect 2494 2347 5434 701997
rect 6214 2347 9154 701997
rect 9934 2347 12874 701997
rect 13654 2347 16594 701997
rect 17374 2347 20314 701997
rect 21094 2347 24034 701997
rect 24814 2347 27754 701997
rect 28534 2347 37714 701997
rect 38494 2347 41434 701997
rect 42214 2347 45154 701997
rect 45934 2347 48874 701997
rect 49654 2347 52594 701997
rect 53374 2347 56314 701997
rect 57094 2347 60034 701997
rect 60814 2347 63754 701997
rect 64534 645876 73714 701997
rect 74494 645876 77434 701997
rect 78214 646060 81154 701997
rect 81934 646060 84874 701997
rect 78214 645876 84874 646060
rect 85654 645876 88594 701997
rect 89374 646060 92314 701997
rect 93094 646060 96034 701997
rect 89374 645876 96034 646060
rect 96814 645876 99754 701997
rect 100534 645876 109714 701997
rect 110494 646060 113434 701997
rect 114214 646060 117154 701997
rect 110494 645876 117154 646060
rect 117934 646060 120874 701997
rect 121654 646060 124594 701997
rect 117934 645876 124594 646060
rect 125374 646060 128314 701997
rect 129094 646060 132034 701997
rect 125374 645876 132034 646060
rect 132814 646060 135754 701997
rect 136534 646060 145714 701997
rect 146494 646060 149434 701997
rect 132814 645876 149434 646060
rect 150214 646060 153154 701997
rect 153934 646060 156874 701997
rect 150214 645876 156874 646060
rect 157654 646060 160594 701997
rect 161374 646060 164314 701997
rect 157654 645876 164314 646060
rect 165094 646060 168034 701997
rect 168814 646060 171754 701997
rect 165094 645876 171754 646060
rect 172534 645876 181714 701997
rect 182494 645876 185434 701997
rect 186214 645876 189154 701997
rect 189934 645876 192874 701997
rect 193654 645876 196594 701997
rect 197374 645876 200314 701997
rect 201094 645876 204034 701997
rect 204814 645876 207754 701997
rect 208534 645876 217714 701997
rect 64534 558816 217714 645876
rect 64534 478978 73714 558816
rect 74494 478978 77434 558816
rect 78214 478978 81154 558816
rect 81934 478978 84874 558816
rect 85654 558632 92314 558816
rect 85654 479162 88594 558632
rect 89374 479162 92314 558632
rect 85654 478978 92314 479162
rect 93094 478978 96034 558816
rect 96814 478978 99754 558816
rect 100534 478978 109714 558816
rect 110494 558632 117154 558816
rect 110494 479162 113434 558632
rect 114214 479162 117154 558632
rect 110494 478978 117154 479162
rect 117934 558632 124594 558816
rect 117934 479162 120874 558632
rect 121654 479162 124594 558632
rect 117934 478978 124594 479162
rect 125374 558632 132034 558816
rect 125374 479162 128314 558632
rect 129094 479162 132034 558632
rect 125374 478978 132034 479162
rect 132814 558632 149434 558816
rect 132814 479162 135754 558632
rect 136534 479162 145714 558632
rect 146494 479162 149434 558632
rect 132814 478978 149434 479162
rect 150214 558632 189154 558816
rect 150214 479162 153154 558632
rect 153934 479162 156874 558632
rect 157654 479162 160594 558632
rect 161374 479162 164314 558632
rect 165094 479162 168034 558632
rect 168814 479162 171754 558632
rect 172534 479162 181714 558632
rect 182494 479162 185434 558632
rect 186214 479162 189154 558632
rect 150214 478978 189154 479162
rect 189934 558632 196594 558816
rect 189934 479162 192874 558632
rect 193654 479162 196594 558632
rect 189934 478978 196594 479162
rect 197374 478978 200314 558816
rect 201094 478978 204034 558816
rect 204814 478978 207754 558816
rect 208534 478978 217714 558816
rect 64534 391918 217714 478978
rect 64534 312084 73714 391918
rect 74494 312084 77434 391918
rect 78214 391734 84874 391918
rect 78214 312268 81154 391734
rect 81934 312268 84874 391734
rect 78214 312084 84874 312268
rect 85654 312084 88594 391918
rect 89374 391734 96034 391918
rect 89374 312268 92314 391734
rect 93094 312268 96034 391734
rect 89374 312084 96034 312268
rect 96814 312084 99754 391918
rect 100534 312084 109714 391918
rect 110494 391734 117154 391918
rect 110494 312268 113434 391734
rect 114214 312268 117154 391734
rect 110494 312084 117154 312268
rect 117934 391734 124594 391918
rect 117934 312268 120874 391734
rect 121654 312268 124594 391734
rect 117934 312084 124594 312268
rect 125374 391734 132034 391918
rect 125374 312268 128314 391734
rect 129094 312268 132034 391734
rect 125374 312084 132034 312268
rect 132814 391734 149434 391918
rect 132814 312268 135754 391734
rect 136534 312268 145714 391734
rect 146494 312268 149434 391734
rect 132814 312084 149434 312268
rect 150214 391734 156874 391918
rect 150214 312268 153154 391734
rect 153934 312268 156874 391734
rect 150214 312084 156874 312268
rect 157654 391734 164314 391918
rect 157654 312268 160594 391734
rect 161374 312268 164314 391734
rect 157654 312084 164314 312268
rect 165094 391734 171754 391918
rect 165094 312268 168034 391734
rect 168814 312268 171754 391734
rect 165094 312084 171754 312268
rect 172534 312084 181714 391918
rect 182494 312084 185434 391918
rect 186214 312084 189154 391918
rect 189934 312084 192874 391918
rect 193654 312084 196594 391918
rect 197374 312084 200314 391918
rect 201094 312084 204034 391918
rect 204814 312084 207754 391918
rect 208534 312084 217714 391918
rect 64534 225024 217714 312084
rect 64534 145184 73714 225024
rect 74494 145184 77434 225024
rect 78214 145184 81154 225024
rect 81934 145184 84874 225024
rect 85654 224840 92314 225024
rect 85654 145368 88594 224840
rect 89374 145368 92314 224840
rect 85654 145184 92314 145368
rect 93094 145184 96034 225024
rect 96814 145184 99754 225024
rect 100534 145184 109714 225024
rect 110494 224840 117154 225024
rect 110494 145368 113434 224840
rect 114214 145368 117154 224840
rect 110494 145184 117154 145368
rect 117934 224840 124594 225024
rect 117934 145368 120874 224840
rect 121654 145368 124594 224840
rect 117934 145184 124594 145368
rect 125374 224840 132034 225024
rect 125374 145368 128314 224840
rect 129094 145368 132034 224840
rect 125374 145184 132034 145368
rect 132814 224840 149434 225024
rect 132814 145368 135754 224840
rect 136534 145368 145714 224840
rect 146494 145368 149434 224840
rect 132814 145184 149434 145368
rect 150214 224840 189154 225024
rect 150214 145368 153154 224840
rect 153934 145368 156874 224840
rect 157654 145368 160594 224840
rect 161374 145368 164314 224840
rect 165094 145368 168034 224840
rect 168814 145368 171754 224840
rect 172534 145368 181714 224840
rect 182494 145368 185434 224840
rect 186214 145368 189154 224840
rect 150214 145184 189154 145368
rect 189934 224840 196594 225024
rect 189934 145368 192874 224840
rect 193654 145368 196594 224840
rect 189934 145184 196594 145368
rect 197374 145184 200314 225024
rect 201094 145184 204034 225024
rect 204814 145184 207754 225024
rect 208534 145184 217714 225024
rect 64534 58166 217714 145184
rect 64534 58124 92314 58166
rect 64534 2347 73714 58124
rect 74494 2347 77434 58124
rect 78214 57940 84874 58124
rect 78214 2347 81154 57940
rect 81934 2347 84874 57940
rect 85654 2347 88594 58124
rect 89374 2347 92314 58124
rect 93094 58124 164314 58166
rect 93094 2347 96034 58124
rect 96814 2347 99754 58124
rect 100534 2347 109714 58124
rect 110494 57940 117154 58124
rect 110494 2347 113434 57940
rect 114214 2347 117154 57940
rect 117934 57940 124594 58124
rect 117934 2347 120874 57940
rect 121654 2347 124594 57940
rect 125374 57940 132034 58124
rect 125374 2347 128314 57940
rect 129094 2347 132034 57940
rect 132814 57940 149434 58124
rect 132814 2347 135754 57940
rect 136534 2347 145714 57940
rect 146494 2347 149434 57940
rect 150214 57940 156874 58124
rect 150214 2347 153154 57940
rect 153934 2347 156874 57940
rect 157654 57940 164314 58124
rect 165094 58124 200314 58166
rect 157654 2347 160594 57940
rect 161374 2347 164314 57940
rect 165094 57940 171754 58124
rect 165094 2347 168034 57940
rect 168814 2347 171754 57940
rect 172534 2347 181714 58124
rect 182494 2347 185434 58124
rect 186214 2347 189154 58124
rect 189934 2347 192874 58124
rect 193654 2347 196594 58124
rect 197374 2347 200314 58124
rect 201094 58124 217714 58166
rect 201094 2347 204034 58124
rect 204814 2347 207754 58124
rect 208534 2347 217714 58124
rect 218494 2347 221434 701997
rect 222214 2347 225154 701997
rect 225934 2347 228874 701997
rect 229654 2347 232594 701997
rect 233374 2347 236314 701997
rect 237094 2347 240034 701997
rect 240814 2347 243754 701997
rect 244534 2347 253714 701997
rect 254494 2347 257434 701997
rect 258214 2347 261154 701997
rect 261934 2347 264874 701997
rect 265654 2347 268594 701997
rect 269374 2347 272314 701997
rect 273094 2347 276034 701997
rect 276814 2347 279754 701997
rect 280534 2347 289714 701997
rect 290494 2347 293434 701997
rect 294214 2347 297154 701997
rect 297934 2347 300874 701997
rect 301654 2347 304594 701997
rect 305374 2347 308314 701997
rect 309094 2347 312034 701997
rect 312814 2347 315754 701997
rect 316534 2347 325714 701997
rect 326494 2347 329434 701997
rect 330214 2347 333154 701997
rect 333934 2347 336874 701997
rect 337654 2347 340594 701997
rect 341374 2347 344314 701997
rect 345094 2347 348034 701997
rect 348814 2347 351754 701997
rect 352534 2347 361714 701997
rect 362494 2347 365434 701997
rect 366214 2347 369154 701997
rect 369934 645876 372874 701997
rect 373654 645876 376594 701997
rect 377374 645876 380314 701997
rect 381094 645876 384034 701997
rect 384814 645876 387754 701997
rect 388534 645876 397714 701997
rect 398494 645876 401434 701997
rect 402214 646060 405154 701997
rect 405934 646060 408874 701997
rect 402214 645876 408874 646060
rect 409654 646060 412594 701997
rect 413374 646060 416314 701997
rect 409654 645876 416314 646060
rect 417094 646060 420034 701997
rect 420814 646060 423754 701997
rect 417094 645876 423754 646060
rect 424534 645876 433714 701997
rect 434494 646060 437434 701997
rect 438214 646060 441154 701997
rect 434494 645876 441154 646060
rect 441934 646060 444874 701997
rect 445654 646060 448594 701997
rect 441934 645876 448594 646060
rect 449374 646060 452314 701997
rect 453094 646060 456034 701997
rect 449374 645876 456034 646060
rect 456814 646060 459754 701997
rect 460534 646060 469714 701997
rect 470494 646060 473434 701997
rect 456814 645876 473434 646060
rect 474214 645876 477154 701997
rect 477934 645876 480874 701997
rect 481654 645876 484594 701997
rect 485374 645876 488314 701997
rect 489094 645876 492034 701997
rect 492814 645876 495754 701997
rect 496534 645876 505714 701997
rect 506494 645876 509434 701997
rect 510214 645876 513154 701997
rect 369934 558816 513154 645876
rect 369934 478978 372874 558816
rect 373654 478978 376594 558816
rect 377374 478978 380314 558816
rect 381094 478978 384034 558816
rect 384814 558632 416314 558816
rect 384814 479162 387754 558632
rect 388534 479162 397714 558632
rect 398494 479162 401434 558632
rect 402214 479162 405154 558632
rect 405934 479162 408874 558632
rect 409654 479162 412594 558632
rect 413374 479162 416314 558632
rect 384814 478978 416314 479162
rect 417094 558632 433714 558816
rect 417094 479162 420034 558632
rect 420814 479162 423754 558632
rect 424534 479162 433714 558632
rect 417094 478978 433714 479162
rect 434494 558632 441154 558816
rect 434494 479162 437434 558632
rect 438214 479162 441154 558632
rect 434494 478978 441154 479162
rect 441934 558632 448594 558816
rect 441934 479162 444874 558632
rect 445654 479162 448594 558632
rect 441934 478978 448594 479162
rect 449374 558632 456034 558816
rect 449374 479162 452314 558632
rect 453094 479162 456034 558632
rect 449374 478978 456034 479162
rect 456814 558632 473434 558816
rect 456814 479162 459754 558632
rect 460534 479162 469714 558632
rect 470494 479162 473434 558632
rect 456814 478978 473434 479162
rect 474214 558632 480874 558816
rect 474214 479162 477154 558632
rect 477934 479162 480874 558632
rect 474214 478978 480874 479162
rect 481654 478978 484594 558816
rect 485374 478978 488314 558816
rect 489094 478978 492034 558816
rect 492814 478978 495754 558816
rect 496534 478978 505714 558816
rect 506494 478978 509434 558816
rect 510214 478978 513154 558816
rect 369934 391918 513154 478978
rect 369934 312084 372874 391918
rect 373654 312084 376594 391918
rect 377374 312084 380314 391918
rect 381094 312084 384034 391918
rect 384814 312084 387754 391918
rect 388534 312084 397714 391918
rect 398494 312084 401434 391918
rect 402214 391734 408874 391918
rect 402214 312268 405154 391734
rect 405934 312268 408874 391734
rect 402214 312084 408874 312268
rect 409654 391734 416314 391918
rect 409654 312268 412594 391734
rect 413374 312268 416314 391734
rect 409654 312084 416314 312268
rect 417094 391734 423754 391918
rect 417094 312268 420034 391734
rect 420814 312268 423754 391734
rect 417094 312084 423754 312268
rect 424534 312084 433714 391918
rect 434494 391734 441154 391918
rect 434494 312268 437434 391734
rect 438214 312268 441154 391734
rect 434494 312084 441154 312268
rect 441934 391734 448594 391918
rect 441934 312268 444874 391734
rect 445654 312268 448594 391734
rect 441934 312084 448594 312268
rect 449374 391734 456034 391918
rect 449374 312268 452314 391734
rect 453094 312268 456034 391734
rect 449374 312084 456034 312268
rect 456814 391734 473434 391918
rect 456814 312268 459754 391734
rect 460534 312268 469714 391734
rect 470494 312268 473434 391734
rect 456814 312084 473434 312268
rect 474214 312084 477154 391918
rect 477934 312084 480874 391918
rect 481654 312084 484594 391918
rect 485374 312084 488314 391918
rect 489094 312084 492034 391918
rect 492814 312084 495754 391918
rect 496534 312084 505714 391918
rect 506494 312084 509434 391918
rect 510214 312084 513154 391918
rect 369934 225024 513154 312084
rect 369934 145184 372874 225024
rect 373654 145184 376594 225024
rect 377374 145184 380314 225024
rect 381094 145184 384034 225024
rect 384814 224840 416314 225024
rect 384814 145368 387754 224840
rect 388534 145368 397714 224840
rect 398494 145368 401434 224840
rect 402214 145368 405154 224840
rect 405934 145368 408874 224840
rect 409654 145368 412594 224840
rect 413374 145368 416314 224840
rect 384814 145184 416314 145368
rect 417094 224840 433714 225024
rect 417094 145368 420034 224840
rect 420814 145368 423754 224840
rect 424534 145368 433714 224840
rect 417094 145184 433714 145368
rect 434494 224840 441154 225024
rect 434494 145368 437434 224840
rect 438214 145368 441154 224840
rect 434494 145184 441154 145368
rect 441934 224840 448594 225024
rect 441934 145368 444874 224840
rect 445654 145368 448594 224840
rect 441934 145184 448594 145368
rect 449374 224840 456034 225024
rect 449374 145368 452314 224840
rect 453094 145368 456034 224840
rect 449374 145184 456034 145368
rect 456814 224840 473434 225024
rect 456814 145368 459754 224840
rect 460534 145368 469714 224840
rect 470494 145368 473434 224840
rect 456814 145184 473434 145368
rect 474214 224840 480874 225024
rect 474214 145368 477154 224840
rect 477934 145368 480874 224840
rect 474214 145184 480874 145368
rect 481654 145184 484594 225024
rect 485374 145184 488314 225024
rect 489094 145184 492034 225024
rect 492814 145184 495754 225024
rect 496534 145184 505714 225024
rect 506494 145184 509434 225024
rect 510214 145184 513154 225024
rect 369934 58166 513154 145184
rect 369934 58124 380314 58166
rect 369934 2347 372874 58124
rect 373654 2347 376594 58124
rect 377374 2347 380314 58124
rect 381094 58124 416314 58166
rect 381094 2347 384034 58124
rect 384814 2347 387754 58124
rect 388534 2347 397714 58124
rect 398494 2347 401434 58124
rect 402214 57940 408874 58124
rect 402214 2347 405154 57940
rect 405934 2347 408874 57940
rect 409654 57940 416314 58124
rect 417094 58124 488314 58166
rect 409654 2347 412594 57940
rect 413374 2347 416314 57940
rect 417094 57940 423754 58124
rect 417094 2347 420034 57940
rect 420814 2347 423754 57940
rect 424534 2347 433714 58124
rect 434494 57940 441154 58124
rect 434494 2347 437434 57940
rect 438214 2347 441154 57940
rect 441934 57940 448594 58124
rect 441934 2347 444874 57940
rect 445654 2347 448594 57940
rect 449374 57940 456034 58124
rect 449374 2347 452314 57940
rect 453094 2347 456034 57940
rect 456814 57940 473434 58124
rect 456814 2347 459754 57940
rect 460534 2347 469714 57940
rect 470494 2347 473434 57940
rect 474214 2347 477154 58124
rect 477934 2347 480874 58124
rect 481654 2347 484594 58124
rect 485374 2347 488314 58124
rect 489094 58124 513154 58166
rect 489094 2347 492034 58124
rect 492814 2347 495754 58124
rect 496534 2347 505714 58124
rect 506494 2347 509434 58124
rect 510214 2347 513154 58124
rect 513934 2347 516874 701997
rect 517654 2347 520594 701997
rect 521374 2347 524314 701997
rect 525094 2347 528034 701997
rect 528814 2347 531754 701997
rect 532534 2347 541714 701997
rect 542494 2347 545434 701997
rect 546214 2347 549154 701997
rect 549934 2347 552874 701997
rect 553654 2347 556594 701997
rect 557374 2347 560314 701997
rect 561094 2347 564034 701997
rect 564814 2347 567754 701997
rect 568534 2347 575309 701997
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 698026 592650 698646
rect -8726 694306 592650 694926
rect -8726 690586 592650 691206
rect -8726 686866 592650 687486
rect -8726 676906 592650 677526
rect -8726 673186 592650 673806
rect -8726 669466 592650 670086
rect -8726 665746 592650 666366
rect -8726 662026 592650 662646
rect -8726 658306 592650 658926
rect -8726 654586 592650 655206
rect -8726 650866 592650 651486
rect -8726 640906 592650 641526
rect -8726 637186 592650 637806
rect -8726 633466 592650 634086
rect -8726 629746 592650 630366
rect -8726 626026 592650 626646
rect -8726 622306 592650 622926
rect -8726 618586 592650 619206
rect -8726 614866 592650 615486
rect -8726 604906 592650 605526
rect -8726 601186 592650 601806
rect -8726 597466 592650 598086
rect -8726 593746 592650 594366
rect -8726 590026 592650 590646
rect -8726 586306 592650 586926
rect -8726 582586 592650 583206
rect -8726 578866 592650 579486
rect -8726 568906 592650 569526
rect -8726 565186 592650 565806
rect -8726 561466 592650 562086
rect -8726 557746 592650 558366
rect -8726 554026 592650 554646
rect -8726 550306 592650 550926
rect -8726 546586 592650 547206
rect -8726 542866 592650 543486
rect -8726 532906 592650 533526
rect -8726 529186 592650 529806
rect -8726 525466 592650 526086
rect -8726 521746 592650 522366
rect -8726 518026 592650 518646
rect -8726 514306 592650 514926
rect -8726 510586 592650 511206
rect -8726 506866 592650 507486
rect -8726 496906 592650 497526
rect -8726 493186 592650 493806
rect -8726 489466 592650 490086
rect -8726 485746 592650 486366
rect -8726 482026 592650 482646
rect -8726 478306 592650 478926
rect -8726 474586 592650 475206
rect -8726 470866 592650 471486
rect -8726 460906 592650 461526
rect -8726 457186 592650 457806
rect -8726 453466 592650 454086
rect -8726 449746 592650 450366
rect -8726 446026 592650 446646
rect -8726 442306 592650 442926
rect -8726 438586 592650 439206
rect -8726 434866 592650 435486
rect -8726 424906 592650 425526
rect -8726 421186 592650 421806
rect -8726 417466 592650 418086
rect -8726 413746 592650 414366
rect -8726 410026 592650 410646
rect -8726 406306 592650 406926
rect -8726 402586 592650 403206
rect -8726 398866 592650 399486
rect -8726 388906 592650 389526
rect -8726 385186 592650 385806
rect -8726 381466 592650 382086
rect -8726 377746 592650 378366
rect -8726 374026 592650 374646
rect -8726 370306 592650 370926
rect -8726 366586 592650 367206
rect -8726 362866 592650 363486
rect -8726 352906 592650 353526
rect -8726 349186 592650 349806
rect -8726 345466 592650 346086
rect -8726 341746 592650 342366
rect -8726 338026 592650 338646
rect -8726 334306 592650 334926
rect -8726 330586 592650 331206
rect -8726 326866 592650 327486
rect -8726 316906 592650 317526
rect -8726 313186 592650 313806
rect -8726 309466 592650 310086
rect -8726 305746 592650 306366
rect -8726 302026 592650 302646
rect -8726 298306 592650 298926
rect -8726 294586 592650 295206
rect -8726 290866 592650 291486
rect -8726 280906 592650 281526
rect -8726 277186 592650 277806
rect -8726 273466 592650 274086
rect -8726 269746 592650 270366
rect -8726 266026 592650 266646
rect -8726 262306 592650 262926
rect -8726 258586 592650 259206
rect -8726 254866 592650 255486
rect -8726 244906 592650 245526
rect -8726 241186 592650 241806
rect -8726 237466 592650 238086
rect -8726 233746 592650 234366
rect -8726 230026 592650 230646
rect -8726 226306 592650 226926
rect -8726 222586 592650 223206
rect -8726 218866 592650 219486
rect -8726 208906 592650 209526
rect -8726 205186 592650 205806
rect -8726 201466 592650 202086
rect -8726 197746 592650 198366
rect -8726 194026 592650 194646
rect -8726 190306 592650 190926
rect -8726 186586 592650 187206
rect -8726 182866 592650 183486
rect -8726 172906 592650 173526
rect -8726 169186 592650 169806
rect -8726 165466 592650 166086
rect -8726 161746 592650 162366
rect -8726 158026 592650 158646
rect -8726 154306 592650 154926
rect -8726 150586 592650 151206
rect -8726 146866 592650 147486
rect -8726 136906 592650 137526
rect -8726 133186 592650 133806
rect -8726 129466 592650 130086
rect -8726 125746 592650 126366
rect -8726 122026 592650 122646
rect -8726 118306 592650 118926
rect -8726 114586 592650 115206
rect -8726 110866 592650 111486
rect -8726 100906 592650 101526
rect -8726 97186 592650 97806
rect -8726 93466 592650 94086
rect -8726 89746 592650 90366
rect -8726 86026 592650 86646
rect -8726 82306 592650 82926
rect -8726 78586 592650 79206
rect -8726 74866 592650 75486
rect -8726 64906 592650 65526
rect -8726 61186 592650 61806
rect -8726 57466 592650 58086
rect -8726 53746 592650 54366
rect -8726 50026 592650 50646
rect -8726 46306 592650 46926
rect -8726 42586 592650 43206
rect -8726 38866 592650 39486
rect -8726 28906 592650 29526
rect -8726 25186 592650 25806
rect -8726 21466 592650 22086
rect -8726 17746 592650 18366
rect -8726 14026 592650 14646
rect -8726 10306 592650 10926
rect -8726 6586 592650 7206
rect -8726 2866 592650 3486
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< obsm5 >>
rect 668 490406 536244 490780
rect 668 486686 536244 489146
rect 668 482966 536244 485426
rect 668 479246 536244 481706
rect 668 475526 536244 477986
rect 668 471806 536244 474266
rect 668 461846 536244 470546
rect 668 458126 536244 460586
rect 668 454406 536244 456866
rect 668 450686 536244 453146
rect 668 446966 536244 449426
rect 668 443246 536244 445706
rect 668 439526 536244 441986
rect 668 435806 536244 438266
rect 668 425846 536244 434546
rect 668 422126 536244 424586
rect 668 418406 536244 420866
rect 668 414686 536244 417146
rect 668 410966 536244 413426
rect 668 407246 536244 409706
rect 668 403526 536244 405986
rect 668 399806 536244 402266
rect 668 389846 536244 398546
rect 668 386126 536244 388586
rect 668 382406 536244 384866
rect 668 378686 536244 381146
rect 668 374966 536244 377426
rect 668 371246 536244 373706
rect 668 367526 536244 369986
rect 668 363806 536244 366266
rect 668 353846 536244 362546
rect 668 350126 536244 352586
rect 668 346406 536244 348866
rect 668 342686 536244 345146
rect 668 338966 536244 341426
rect 668 335246 536244 337706
rect 668 331526 536244 333986
rect 668 327806 536244 330266
rect 668 317846 536244 326546
rect 668 314126 536244 316586
rect 668 310406 536244 312866
rect 668 306686 536244 309146
rect 668 302966 536244 305426
rect 668 299246 536244 301706
rect 668 295526 536244 297986
rect 668 291806 536244 294266
rect 668 281846 536244 290546
rect 668 278126 536244 280586
rect 668 274406 536244 276866
rect 668 270686 536244 273146
rect 668 266966 536244 269426
rect 668 263246 536244 265706
rect 668 259526 536244 261986
rect 668 255806 536244 258266
rect 668 245846 536244 254546
rect 668 242126 536244 244586
rect 668 238406 536244 240866
rect 668 234686 536244 237146
rect 668 230966 536244 233426
rect 668 227246 536244 229706
rect 668 223526 536244 225986
rect 668 219806 536244 222266
rect 668 209846 536244 218546
rect 668 206126 536244 208586
rect 668 202406 536244 204866
rect 668 198686 536244 201146
rect 668 194966 536244 197426
rect 668 191246 536244 193706
rect 668 187526 536244 189986
rect 668 183806 536244 186266
rect 668 173846 536244 182546
rect 668 170126 536244 172586
rect 668 166406 536244 168866
rect 668 162686 536244 165146
rect 668 158966 536244 161426
rect 668 155246 536244 157706
rect 668 151526 536244 153986
rect 668 147806 536244 150266
rect 668 145700 536244 146546
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 1794 -7654 2414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 -7654 38414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 -7654 74414 58044 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 145264 74414 224944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 312164 74414 391838 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 479058 74414 558736 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 645956 74414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 -7654 110414 58044 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 145264 110414 224944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 312164 110414 391838 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 479058 110414 558736 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 645956 110414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 -7654 146414 57860 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 145448 146414 224760 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 312348 146414 391654 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 479242 146414 558552 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 646140 146414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 -7654 182414 58044 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 145448 182414 224760 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 312164 182414 391838 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 479242 182414 558552 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 645956 182414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 -7654 218414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 -7654 254414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 -7654 290414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 -7654 326414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 -7654 362414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 -7654 398414 58044 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 145448 398414 224760 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 312164 398414 391838 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 479242 398414 558552 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 645956 398414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 -7654 434414 58044 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 145264 434414 224944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 312164 434414 391838 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 479058 434414 558736 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 645956 434414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 -7654 470414 57860 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 145448 470414 224760 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 312348 470414 391654 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 479242 470414 558552 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 646140 470414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 -7654 506414 58044 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 145264 506414 224944 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 312164 506414 391838 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 479058 506414 558736 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 645956 506414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 -7654 542414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 577794 -7654 578414 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 2866 592650 3486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 38866 592650 39486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 74866 592650 75486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 110866 592650 111486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 146866 592650 147486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 182866 592650 183486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 218866 592650 219486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 254866 592650 255486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 290866 592650 291486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 326866 592650 327486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 362866 592650 363486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 398866 592650 399486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 434866 592650 435486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 470866 592650 471486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 506866 592650 507486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 542866 592650 543486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 578866 592650 579486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 614866 592650 615486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 650866 592650 651486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 686866 592650 687486 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 9234 -7654 9854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 45234 -7654 45854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 81234 -7654 81854 57860 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 81234 145264 81854 224944 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 81234 312348 81854 391654 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 81234 479058 81854 558736 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 81234 646140 81854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 117234 -7654 117854 58044 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 117234 145264 117854 224944 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 117234 312164 117854 391838 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 117234 479058 117854 558736 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 117234 645956 117854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 153234 -7654 153854 57860 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 153234 145448 153854 224760 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 153234 312348 153854 391654 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 153234 479242 153854 558552 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 153234 646140 153854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 189234 -7654 189854 58044 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 189234 145264 189854 224944 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 189234 312164 189854 391838 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 189234 479058 189854 558736 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 189234 645956 189854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 225234 -7654 225854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 261234 -7654 261854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 297234 -7654 297854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 333234 -7654 333854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 369234 -7654 369854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 405234 -7654 405854 57860 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 405234 145448 405854 224760 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 405234 312348 405854 391654 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 405234 479242 405854 558552 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 405234 646140 405854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 441234 -7654 441854 58044 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 441234 145264 441854 224944 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 441234 312164 441854 391838 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 441234 479058 441854 558736 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 441234 645956 441854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 477234 -7654 477854 58044 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 477234 145448 477854 224760 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 477234 312164 477854 391838 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 477234 479242 477854 558552 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 477234 645956 477854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 513234 -7654 513854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 549234 -7654 549854 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 10306 592650 10926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 46306 592650 46926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 82306 592650 82926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 118306 592650 118926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 154306 592650 154926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 190306 592650 190926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 226306 592650 226926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 262306 592650 262926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 298306 592650 298926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 334306 592650 334926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 370306 592650 370926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 406306 592650 406926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 442306 592650 442926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 478306 592650 478926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 514306 592650 514926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 550306 592650 550926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 586306 592650 586926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 622306 592650 622926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 658306 592650 658926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 694306 592650 694926 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 16674 -7654 17294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 52674 -7654 53294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 88674 -7654 89294 58044 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 88674 145448 89294 224760 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 88674 312164 89294 391838 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 88674 479242 89294 558552 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 88674 645956 89294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 124674 -7654 125294 58044 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 124674 145264 125294 224944 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 124674 312164 125294 391838 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 124674 479058 125294 558736 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 124674 645956 125294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 160674 -7654 161294 57860 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 160674 145448 161294 224760 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 160674 312348 161294 391654 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 160674 479242 161294 558552 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 160674 646140 161294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 196674 -7654 197294 58044 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 196674 145264 197294 224944 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 196674 312164 197294 391838 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 196674 479058 197294 558736 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 196674 645956 197294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 232674 -7654 233294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 268674 -7654 269294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 304674 -7654 305294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 340674 -7654 341294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 376674 -7654 377294 58044 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 376674 145264 377294 224944 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 376674 312164 377294 391838 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 376674 479058 377294 558736 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 376674 645956 377294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 412674 -7654 413294 57860 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 412674 145448 413294 224760 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 412674 312348 413294 391654 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 412674 479242 413294 558552 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 412674 646140 413294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 448674 -7654 449294 58044 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 448674 145264 449294 224944 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 448674 312164 449294 391838 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 448674 479058 449294 558736 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 448674 645956 449294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 484674 -7654 485294 58044 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 484674 145264 485294 224944 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 484674 312164 485294 391838 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 484674 479058 485294 558736 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 484674 645956 485294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 520674 -7654 521294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 556674 -7654 557294 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 17746 592650 18366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 53746 592650 54366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 89746 592650 90366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 125746 592650 126366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 161746 592650 162366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 197746 592650 198366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 233746 592650 234366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 269746 592650 270366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 305746 592650 306366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 341746 592650 342366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 377746 592650 378366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 413746 592650 414366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 449746 592650 450366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 485746 592650 486366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 521746 592650 522366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 557746 592650 558366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 593746 592650 594366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 629746 592650 630366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 665746 592650 666366 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 24114 -7654 24734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 60114 -7654 60734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 96114 -7654 96734 58044 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 96114 145264 96734 224944 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 96114 312164 96734 391838 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 96114 479058 96734 558736 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 96114 645956 96734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 132114 -7654 132734 58044 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 132114 145264 132734 224944 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 132114 312164 132734 391838 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 132114 479058 132734 558736 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 132114 645956 132734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 168114 -7654 168734 57860 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 168114 145448 168734 224760 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 168114 312348 168734 391654 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 168114 479242 168734 558552 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 168114 646140 168734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 204114 -7654 204734 58044 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 204114 145264 204734 224944 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 204114 312164 204734 391838 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 204114 479058 204734 558736 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 204114 645956 204734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 240114 -7654 240734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 276114 -7654 276734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 312114 -7654 312734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 348114 -7654 348734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 384114 -7654 384734 58044 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 384114 145264 384734 224944 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 384114 312164 384734 391838 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 384114 479058 384734 558736 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 384114 645956 384734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 420114 -7654 420734 57860 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 420114 145448 420734 224760 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 420114 312348 420734 391654 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 420114 479242 420734 558552 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 420114 646140 420734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 456114 -7654 456734 58044 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 456114 145264 456734 224944 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 456114 312164 456734 391838 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 456114 479058 456734 558736 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 456114 645956 456734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 492114 -7654 492734 58044 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 492114 145264 492734 224944 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 492114 312164 492734 391838 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 492114 479058 492734 558736 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 492114 645956 492734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 528114 -7654 528734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 564114 -7654 564734 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 25186 592650 25806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 61186 592650 61806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 97186 592650 97806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 133186 592650 133806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 169186 592650 169806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 205186 592650 205806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 241186 592650 241806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 277186 592650 277806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 313186 592650 313806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 349186 592650 349806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 385186 592650 385806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 421186 592650 421806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 457186 592650 457806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 493186 592650 493806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 529186 592650 529806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 565186 592650 565806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 601186 592650 601806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 637186 592650 637806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 673186 592650 673806 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 20394 -7654 21014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 56394 -7654 57014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 92394 -7654 93014 58086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 92394 145264 93014 224944 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 92394 312348 93014 391654 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 92394 479058 93014 558736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 92394 646140 93014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 128394 -7654 129014 57860 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 128394 145448 129014 224760 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 128394 312348 129014 391654 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 128394 479242 129014 558552 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 128394 646140 129014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 164394 -7654 165014 58086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 164394 145448 165014 224760 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 164394 312164 165014 391838 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 164394 479242 165014 558552 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 164394 645956 165014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 200394 -7654 201014 58086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 200394 145264 201014 224944 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 200394 312164 201014 391838 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 200394 479058 201014 558736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 200394 645956 201014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 236394 -7654 237014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 272394 -7654 273014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 308394 -7654 309014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 344394 -7654 345014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 380394 -7654 381014 58086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 380394 145264 381014 224944 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 380394 312164 381014 391838 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 380394 479058 381014 558736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 380394 645956 381014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 416394 -7654 417014 58086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 416394 145264 417014 224944 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 416394 312164 417014 391838 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 416394 479058 417014 558736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 416394 645956 417014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 452394 -7654 453014 57860 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 452394 145448 453014 224760 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 452394 312348 453014 391654 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 452394 479242 453014 558552 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 452394 646140 453014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 488394 -7654 489014 58086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 488394 145264 489014 224944 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 488394 312164 489014 391838 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 488394 479058 489014 558736 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 488394 645956 489014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 524394 -7654 525014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 560394 -7654 561014 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 21466 592650 22086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 57466 592650 58086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 93466 592650 94086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 129466 592650 130086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 165466 592650 166086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 201466 592650 202086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 237466 592650 238086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 273466 592650 274086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 309466 592650 310086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 345466 592650 346086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 381466 592650 382086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 417466 592650 418086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 453466 592650 454086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 489466 592650 490086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 525466 592650 526086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 561466 592650 562086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 597466 592650 598086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 633466 592650 634086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 669466 592650 670086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 27834 -7654 28454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 63834 -7654 64454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 99834 -7654 100454 58044 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 99834 145264 100454 224944 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 99834 312164 100454 391838 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 99834 479058 100454 558736 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 99834 645956 100454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 135834 -7654 136454 57860 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 135834 145448 136454 224760 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 135834 312348 136454 391654 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 135834 479242 136454 558552 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 135834 646140 136454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 171834 -7654 172454 58044 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 171834 145448 172454 224760 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 171834 312164 172454 391838 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 171834 479242 172454 558552 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 171834 645956 172454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 207834 -7654 208454 58044 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 207834 145264 208454 224944 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 207834 312164 208454 391838 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 207834 479058 208454 558736 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 207834 645956 208454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 243834 -7654 244454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 279834 -7654 280454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 315834 -7654 316454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 351834 -7654 352454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 387834 -7654 388454 58044 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 387834 145448 388454 224760 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 387834 312164 388454 391838 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 387834 479242 388454 558552 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 387834 645956 388454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 423834 -7654 424454 58044 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 423834 145448 424454 224760 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 423834 312164 424454 391838 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 423834 479242 424454 558552 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 423834 645956 424454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 459834 -7654 460454 57860 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 459834 145448 460454 224760 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 459834 312348 460454 391654 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 459834 479242 460454 558552 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 459834 646140 460454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 495834 -7654 496454 58044 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 495834 145264 496454 224944 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 495834 312164 496454 391838 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 495834 479058 496454 558736 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 495834 645956 496454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 531834 -7654 532454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 567834 -7654 568454 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 28906 592650 29526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 64906 592650 65526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 100906 592650 101526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 136906 592650 137526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 172906 592650 173526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 208906 592650 209526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 244906 592650 245526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 280906 592650 281526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 316906 592650 317526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 352906 592650 353526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 388906 592650 389526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 424906 592650 425526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 460906 592650 461526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 496906 592650 497526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 532906 592650 533526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 568906 592650 569526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 604906 592650 605526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 640906 592650 641526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 676906 592650 677526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 5514 -7654 6134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 41514 -7654 42134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 -7654 78134 58044 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 145264 78134 224944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 312164 78134 391838 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 479058 78134 558736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 645956 78134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 -7654 114134 57860 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 145448 114134 224760 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 312348 114134 391654 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 479242 114134 558552 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 646140 114134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149514 -7654 150134 58044 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149514 145264 150134 224944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149514 312164 150134 391838 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149514 479058 150134 558736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149514 645956 150134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 185514 -7654 186134 58044 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 185514 145448 186134 224760 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 185514 312164 186134 391838 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 185514 479242 186134 558552 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 185514 645956 186134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 221514 -7654 222134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 257514 -7654 258134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 293514 -7654 294134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 329514 -7654 330134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 365514 -7654 366134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 -7654 402134 58044 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 145448 402134 224760 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 312164 402134 391838 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 479242 402134 558552 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 645956 402134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 -7654 438134 57860 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 145448 438134 224760 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 312348 438134 391654 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 479242 438134 558552 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 646140 438134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 473514 -7654 474134 58044 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 473514 145264 474134 224944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 473514 312164 474134 391838 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 473514 479058 474134 558736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 473514 645956 474134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 509514 -7654 510134 58044 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 509514 145264 510134 224944 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 509514 312164 510134 391838 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 509514 479058 510134 558736 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 509514 645956 510134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 545514 -7654 546134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 581514 -7654 582134 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 6586 592650 7206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 42586 592650 43206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 78586 592650 79206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 114586 592650 115206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 150586 592650 151206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 186586 592650 187206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 222586 592650 223206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 258586 592650 259206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 294586 592650 295206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 330586 592650 331206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 366586 592650 367206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 402586 592650 403206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 438586 592650 439206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 474586 592650 475206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 510586 592650 511206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 546586 592650 547206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 582586 592650 583206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 618586 592650 619206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 654586 592650 655206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 690586 592650 691206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 12954 -7654 13574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 48954 -7654 49574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 84954 -7654 85574 58044 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 84954 145264 85574 224944 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 84954 312164 85574 391838 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 84954 479058 85574 558736 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 84954 645956 85574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 120954 -7654 121574 57860 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 120954 145448 121574 224760 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 120954 312348 121574 391654 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 120954 479242 121574 558552 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 120954 646140 121574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 156954 -7654 157574 58044 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 156954 145448 157574 224760 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 156954 312164 157574 391838 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 156954 479242 157574 558552 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 156954 645956 157574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192954 -7654 193574 58044 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192954 145448 193574 224760 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192954 312164 193574 391838 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192954 479242 193574 558552 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192954 645956 193574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 228954 -7654 229574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 264954 -7654 265574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 300954 -7654 301574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 336954 -7654 337574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 -7654 373574 58044 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 145264 373574 224944 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 312164 373574 391838 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 479058 373574 558736 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 645956 373574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 408954 -7654 409574 58044 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 408954 145448 409574 224760 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 408954 312164 409574 391838 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 408954 479242 409574 558552 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 408954 645956 409574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444954 -7654 445574 57860 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444954 145448 445574 224760 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444954 312348 445574 391654 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444954 479242 445574 558552 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444954 646140 445574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 480954 -7654 481574 58044 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 480954 145264 481574 224944 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 480954 312164 481574 391838 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 480954 479058 481574 558736 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 480954 645956 481574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 516954 -7654 517574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 552954 -7654 553574 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 14026 592650 14646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 50026 592650 50646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 86026 592650 86646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 122026 592650 122646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 158026 592650 158646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 194026 592650 194646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 230026 592650 230646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 266026 592650 266646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 302026 592650 302646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 338026 592650 338646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 374026 592650 374646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 410026 592650 410646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 446026 592650 446646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 482026 592650 482646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 518026 592650 518646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 554026 592650 554646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 590026 592650 590646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 626026 592650 626646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 662026 592650 662646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 698026 592650 698646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 311604168
string GDS_FILE /home/prherrma/runners/r1/_work/tapeout-ci-2311/tapeout-ci-2311/openlane/user_project_wrapper/runs/23_11_05_22_06/results/signoff/user_project_wrapper.magic.gds
string GDS_START 17101132
<< end >>

