`ifndef CLAM_DEFS_SVH
`define CLAM_DEFS_SVH

/////////////////////////
// BOOT SELECT DEFINES //
/////////////////////////

`define BOOT_NORMAL 0
`define BOOT_FAILSAFE 1

/////////////////////////
// PERIPHERAL DEFINES  //
/////////////////////////

`define SOC_NUM_INTER       54
// `include "Peripheral_Unit_Defs"

`endif // CLAM_DEFS_SVH
