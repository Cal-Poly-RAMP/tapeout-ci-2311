`timescale 1ns / 1ps

///////////////////////////////////////////////////////////////////////////////
//
// Module Name: SPI_Master
// Description: SPI (Serial Peripheral Interface) Master
//              Creates master based on input configuration.
//              Sends a byte one bit at a time on MOSI
//              Will also receive byte data one bit at a time on MISO.
//              Any data on input byte will be shipped out on MOSI.
//
//              To kick-off transaction, user must pulse i_TX_DV.
//              This module supports multi-byte transmissions by pulsing
//              i_TX_DV and loading up i_TX_Byte when o_TX_Ready is high.
//
//              This module is only responsible for controlling Clk, MOSI, 
//              and MISO.  If the SPI peripheral requires a chip-select, 
//              this must be done at a higher level.
//
// Note:        i_Clk must be at least 2x faster than i_SPI_Clk
//
// Config:      i_spi_mode, can be 0, 1, 2, or 3.  See above.
//              Can be configured in one of 4 modes:
//              Mode | Clock Polarity (CPOL/CKP) | Clock Phase (CPHA)
//               0   |             0             |        0
//               1   |             0             |        1
//               2   |             1             |        0
//               3   |             1             |        1
//              More: https://en.wikipedia.org/wiki/Serial_Peripheral_Interface_Bus#Mode_numbers
//              i_ticks_per_half_bit - Sets frequency of o_SPI_Clk.  o_SPI_Clk is
//              derived from i_Clk.  Set to integer number of clocks for each
//              half-bit of SPI data.  E.g. 100 MHz i_Clk, CLKS_PER_HALF_BIT = 2
//              would create o_SPI_CLK of 25 MHz.  Must be >= 2
//
// SPDX-License-Identifier: Apache-2.0
//
///////////////////////////////////////////////////////////////////////////////

module SPI_Master (
   // Control/Data Signals,
   input        i_Rst_L,     // FPGA Reset
   input        i_Clk,       // FPGA Clock
   input        i_wr_cr,
   input        i_wr_data,
   input [1:0]  i_spi_mode,
   input [15:0] i_ticks_per_half_bit,
   input [3:0]  i_data_length,    // Length of data to be transmitted/received minus 1
   
   // TX (MOSI) Signals
   input [15:0] i_TX_Data,        // Data to transmit on MOSI
   input        i_TX_MSB_first,   // Data sent MSB first
   input        i_TX_DV,          // Data Valid Pulse with i_TX_Byte
   output reg   o_TX_Ready,       // Transmit Ready for next byte
   
   // RX (MISO) Signals
   input        i_RX_MSB_first,  // Data received MSB first
   output reg       o_RX_DV,     // Data Valid pulse (1 clock cycle)
   output reg [15:0] o_RX_Data,   // Data received on MISO

   // SPI Interface
   output reg o_SPI_Clk,
   input      i_SPI_MISO,
   output reg o_SPI_MOSI
   );

  // SPI Interface (All Runs at SPI Clock Domain)
  wire w_CPOL;     // Clock polarity
  wire w_CPHA;     // Clock phase

  logic r1_wr_cr = 0, r2_wr_cr = 0, wr_cr;
  logic r1_wr_data = 0, r2_wr_data = 0, wr_data;
  logic [1:0] r_spi_mode = 2'b0;
  logic [15:0] r_ticks_per_half_bit;
  logic [15:0] r_SPI_Clk_Count;
  logic r_SPI_Clk;
  logic [5:0] r_SPI_Clk_Edges;
  logic r_Leading_Edge;
  logic r_Trailing_Edge;
  logic       r_TX_DV;
  logic [3:0] r_data_length;
  logic [5:0] r_data_length_sig;
  logic r_TX_MSB_first;
  logic r_RX_MSB_first;
  logic [15:0] r_TX_Data;

  logic [3:0] r_RX_Bit_Count;
  logic [3:0] r_TX_Bit_Count;

  // CPOL: Clock Polarity
  // CPOL=0 means clock idles at 0, leading edge is rising edge.
  // CPOL=1 means clock idles at 1, leading edge is falling edge.
  assign w_CPOL  = (r_spi_mode == 2) | (r_spi_mode == 3);

  // CPHA: Clock Phase
  // CPHA=0 means the "out" side changes the data on trailing edge of clock
  //              the "in" side captures data on leading edge of clock
  // CPHA=1 means the "out" side changes the data on leading edge of clock
  //              the "in" side captures data on the trailing edge of clock
  assign w_CPHA  = (r_spi_mode == 1) | (r_spi_mode == 3);

  assign wr_cr = r1_wr_cr & ~r2_wr_cr;
  assign wr_data = r1_wr_data & ~r2_wr_data;
  
  assign r_data_length_sig = {2'b0, r_data_length};

  // Purpose: Generate SPI Clock correct number of times when DV pulse comes
  always @(posedge i_Clk)
  begin
    if (~i_Rst_L)
    begin
      o_TX_Ready      <= 1'b0;
      r_spi_mode      <= 0;
      r_ticks_per_half_bit <= 0;
      r_SPI_Clk_Edges <= 0;
      r_TX_MSB_first  <= 0;
      r_RX_MSB_first  <= 0;
      r_Leading_Edge  <= 1'b0;
      r_Trailing_Edge <= 1'b0;
      r_SPI_Clk       <= w_CPOL; // assign default state to idle state
      r_SPI_Clk_Count <= 0;
    end
    else
    begin

      // Default assignments
      r_Leading_Edge  <= 1'b0;
      r_Trailing_Edge <= 1'b0;
      r1_wr_cr <= i_wr_cr;
      r2_wr_cr <= r1_wr_cr;
      r1_wr_data <= i_wr_data;
      r2_wr_data <= r1_wr_data;
      if (wr_cr) begin
          r_spi_mode      <= i_spi_mode;
          r_ticks_per_half_bit <= i_ticks_per_half_bit;
          r_data_length <= i_data_length;
          r_TX_MSB_first <= i_TX_MSB_first;
          r_RX_MSB_first <= i_RX_MSB_first;
      end
      
      if (i_TX_DV)
      begin
        o_TX_Ready      <= 1'b0;
        r_SPI_Clk_Edges <= (r_data_length_sig + 1) << 1;  // Total # edges in data is 2 * (i_TX_data_length + 1)
      end
      else if (r_SPI_Clk_Edges > 0)
      begin
        o_TX_Ready <= 1'b0;
        
        if (r_SPI_Clk_Count == r_ticks_per_half_bit*2-1)
        begin
          r_SPI_Clk_Edges <= r_SPI_Clk_Edges - 1'b1;
          r_Trailing_Edge <= 1'b1;
          r_SPI_Clk_Count <= 0;
          r_SPI_Clk       <= ~r_SPI_Clk;
        end
        else if (r_SPI_Clk_Count == r_ticks_per_half_bit-1)
        begin
          r_SPI_Clk_Edges <= r_SPI_Clk_Edges - 1'b1;
          r_Leading_Edge  <= 1'b1;
          r_SPI_Clk_Count <= r_SPI_Clk_Count + 1'b1;
          r_SPI_Clk       <= ~r_SPI_Clk;
        end
        else
        begin
          r_SPI_Clk_Count <= r_SPI_Clk_Count + 1'b1;
        end
      end  
      else
      begin
        o_TX_Ready <= 1'b1;
      end
      
      
    end // else: !if(~i_Rst_L)
  end // always @ (posedge i_Clk)


  // Purpose: Register i_TX_Byte when Data Valid is pulsed.
  // Keeps local storage of byte in case higher level module changes the data
  always @(posedge i_Clk)
  begin
    if (~i_Rst_L)
    begin
      r_TX_Data <= 16'h0;
      r_TX_DV   <= 1'b0;
    end
    else
      begin
        r_TX_DV <= i_TX_DV; // 1 clock cycle delay
        if (wr_data)
        begin
          r_TX_Data <= i_TX_Data;
        end
      end // else: !if(~i_Rst_L)
  end // always @ (posedge i_Clk)


  // Purpose: Generate MOSI data
  // Works with both CPHA=0 and CPHA=1
  always @(posedge i_Clk)
  begin
    if (~i_Rst_L)
    begin
      o_SPI_MOSI     <= 1'b0;
      r_TX_Bit_Count <= 4'b1111; // send MSb first
    end
    else
    begin
      // If ready is high, reset bit counts to default
      if (o_TX_Ready)
      begin
        if (r_TX_MSB_first)
          r_TX_Bit_Count <= r_data_length;
        else
          r_TX_Bit_Count <= 4'b0;
      end
      // Catch the case where we start transaction and CPHA = 0
      else if (r_TX_DV & ~w_CPHA)
      begin
        if (r_TX_MSB_first) begin
          o_SPI_MOSI     <= r_TX_Data[r_data_length];
          r_TX_Bit_Count <= r_data_length - 1;
        end
        else begin
          o_SPI_MOSI     <= r_TX_Data[0];
          r_TX_Bit_Count <= 4'd1;
        end
      end
      else if ((r_Leading_Edge & w_CPHA) | (r_Trailing_Edge & ~w_CPHA))
      begin
        if (r_TX_MSB_first)
          r_TX_Bit_Count <= r_TX_Bit_Count - 1'b1;
        else
          r_TX_Bit_Count <= r_TX_Bit_Count + 1'b1;
        o_SPI_MOSI     <= r_TX_Data[r_TX_Bit_Count];
      end
    end
  end


  // Purpose: Read in MISO data.
  always @(posedge i_Clk)
  begin
    if (~i_Rst_L)
    begin
      o_RX_Data      <= 16'h0;
      o_RX_DV        <= 1'b0;
      r_RX_Bit_Count <= 4'b1111;
    end
    else
    begin

      // Default Assignments
      o_RX_DV   <= 1'b0;

      if (o_TX_Ready) // Check if ready is high, if so reset bit count to default
      begin
        if (r_RX_MSB_first)
          r_RX_Bit_Count <= r_data_length;
        else
          r_RX_Bit_Count <= 4'b0;
      end
      else if ((r_Leading_Edge & ~w_CPHA) | (r_Trailing_Edge & w_CPHA))
      begin
        if (r_RX_MSB_first)
          r_RX_Bit_Count <= r_RX_Bit_Count - 1'b1;
        else
          r_RX_Bit_Count <= r_RX_Bit_Count + 1'b1;
        o_RX_Data[r_RX_Bit_Count] <= i_SPI_MISO;  // Sample data
        if (r_RX_MSB_first) begin
          if (r_RX_Bit_Count == 4'b0000)
          begin
            o_RX_DV   <= 1'b1;   // Byte done, pulse Data Valid
          end
        end
        else begin
          if (r_RX_Bit_Count == r_data_length)
          begin
            o_RX_DV   <= 1'b1;   // Byte done, pulse Data Valid
          end
        end
      end
    end
  end
  
  
  // Purpose: Add clock delay to signals for alignment.
  always @(posedge i_Clk)
  begin
    if (~i_Rst_L)
    begin
      o_SPI_Clk  <= w_CPOL;
    end
    else
      begin
        o_SPI_Clk <= r_SPI_Clk;
      end // else: !if(~i_Rst_L)
  end // always @ (posedge i_Clk)
  

endmodule // SPI_Master
